package pkg;
        `include "define.svh"
        `include "transaction.sv"
        `include "generator.sv"
        `include "driver.sv"
        `include "reference.sv"
        `include "monitor.sv"
        `include "scoreboard.sv"
        `include "environment.sv"
        `include "test.sv"
endpackage
