parameter W = 8;
parameter num = 10;
parameter SHIFT_WIDTH = $clog2(W);
